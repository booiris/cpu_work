`timescale 1ns / 1ps
`include "defines.v"

module ex(

    );
endmodule
