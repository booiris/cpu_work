`timescale 1ns / 1ps
`include "defines.v"

// 本模块为译码过程

module id(
        input wire rst,
        input wire[`inst_addr_bus] inst_addr,
        input wire[`inst_bus] inst

        
    );
endmodule
