`timescale 1ns / 1ps
`include "defines.v"

// 本模块为译码转向执行的过程


module id_to_ex(

    );
endmodule
