`timescale 1ns / 1ps
`include "defines.v"

// 本模块为 mips 中 32个寄存器的实现

module reg_build(
    
    );
endmodule
